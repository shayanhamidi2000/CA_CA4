module HazardUnit();

endmodule
